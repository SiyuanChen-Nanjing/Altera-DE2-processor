`timescale 1 ns / 100 ps

module processor_tb();

	
	reg clock, reset;
	wire [31:0] alu_result, data_writeReg, data_readRegA, data_readRegB, 
	imm_sx, inst_exec, q_imem, alu_data_inA, alu_data_inB;
	wire [11:0] address_imem;
	wire ctrl_writeEnable;
	wire [4:0] ctrl_writeReg;

	skeleton sk(clock, reset);
	
	initial
	
		begin
			clock = 1'b0;
			reset = 1'b1;
			@(posedge clock);
			reset = 1'b0;
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			@(posedge clock);
			$display("address_imem: %d", address_imem);
			$display("alu_result: %b", alu_result);
			$display("alu_data_inA: %b, alu_data_inB: %b", alu_data_inA, alu_data_inB);
			$display("rd: %b", data_writeReg);
			$display("ctrl_writeReg: %b, ctrl_writeEnable: %b", ctrl_writeReg, ctrl_writeEnable);
			@(negedge clock);
			$display("q_imem: %b", q_imem);
			$stop;
		end
	
	always 
		#10 clock = ~clock;

endmodule